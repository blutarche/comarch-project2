module processor( clock,
reset,
serial_in, serial_valid_in, serial_ready_in, serial_rden_out, serial_out,s serial_wren_out
);