module adder(
    input   [31:0]  i,
    output  [31:0]  o
    );
    assign o = i+4;
endmodule